module patgen(
	input pclk,
	output [7:0] sample_out
);

assign sample_out = 8'd0;

endmodule
